`include "key.sv"