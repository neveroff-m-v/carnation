`include "sensor\.sv"