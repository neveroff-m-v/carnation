`include "tactile\.sv"